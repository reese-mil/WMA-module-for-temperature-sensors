`timescale 1ns/1ps

//WMA Calculator Main Module

//Authors: Kate Bailey, Reese Milhone


module main;
    tb_WMA_Calculator tb(); // instantiate the testbench
endmodule

